* Bruce MacKinnon 7-June-2024
*
* A simplistic model of a 1 MHz crystal using an LC series circuit
* NOTE: Need to add Q factor, etc.
.SUBCKT CRYSTAL_1MC a b 
l1 a c 165u
c1 c b 150p
.ENDS



