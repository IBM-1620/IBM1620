* XXX
* 
* https://static.righto.com/sms/XXX.html
* SPICE model of IBM SMS logic card
* Bruce MacKinnon 7-June-2024

.SUBCKT SMS_CARD_XXX a b c d e f g h j k l m n p q r

* Standard aliases for power/ground pins
Rx0 vp12 n 0
Rx1 vn12 m 0
Rx2 gnd j 0 

* PNP transistor:
* Qx nc nb ne mname 

.ENDS


