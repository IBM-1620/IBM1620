* HIZ
* SPICE model of IBM SMS logic card
* Bruce MacKinnon 7-June-2024

.SUBCKT SMS_CARD_HIZ a

r1 a 0 100MEG

.ENDS


