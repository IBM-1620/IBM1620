module sms_card_cd()
